-- Copyright (C) 2016  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition"
-- CREATED		"Thu Mar 19 22:32:33 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY p1 IS 
	PORT
	(
		P0 :  IN  STD_LOGIC;
		P1 :  IN  STD_LOGIC;
		P2 :  IN  STD_LOGIC;
		P3 :  IN  STD_LOGIC;
		P4 :  IN  STD_LOGIC;
		P5 :  IN  STD_LOGIC;
		P6 :  IN  STD_LOGIC;
		P7 :  IN  STD_LOGIC;
		MR :  IN  STD_LOGIC;
		clock :  IN  STD_LOGIC;
		PSN :  IN  STD_LOGIC;
		LRN :  IN  STD_LOGIC;
		SERIAL :  IN  STD_LOGIC;
		Q0 :  OUT  STD_LOGIC;
		Q1 :  OUT  STD_LOGIC;
		Q2 :  OUT  STD_LOGIC;
		Q3 :  OUT  STD_LOGIC;
		Q4 :  OUT  STD_LOGIC;
		Q5 :  OUT  STD_LOGIC;
		Q6 :  OUT  STD_LOGIC;
		Q7 :  OUT  STD_LOGIC
	);
END p1;

ARCHITECTURE bdf_type OF p1 IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT \74157_0\
	PORT(A1 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 SEL : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 GN : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 Y2 : OUT STD_LOGIC;
		 Y1 : OUT STD_LOGIC;
		 Y4 : OUT STD_LOGIC;
		 Y3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74157_0\: COMPONENT IS true;
ATTRIBUTE noopt OF \74157_0\: COMPONENT IS true;

COMPONENT \74157_3\
	PORT(A1 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 SEL : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 GN : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 Y2 : OUT STD_LOGIC;
		 Y1 : OUT STD_LOGIC;
		 Y4 : OUT STD_LOGIC;
		 Y3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74157_3\: COMPONENT IS true;
ATTRIBUTE noopt OF \74157_3\: COMPONENT IS true;

COMPONENT \74195_1\
	PORT(ST/LDN : IN STD_LOGIC;
		 KN : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 J : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q0 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74195_1\: COMPONENT IS true;
ATTRIBUTE noopt OF \74195_1\: COMPONENT IS true;

COMPONENT \74195_2\
	PORT(ST/LDN : IN STD_LOGIC;
		 KN : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 J : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q0 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74195_2\: COMPONENT IS true;
ATTRIBUTE noopt OF \74195_2\: COMPONENT IS true;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;


BEGIN 
Q0 <= SYNTHESIZED_WIRE_23;
Q1 <= SYNTHESIZED_WIRE_0;
Q2 <= SYNTHESIZED_WIRE_2;
Q3 <= SYNTHESIZED_WIRE_26;
Q4 <= SYNTHESIZED_WIRE_4;
Q5 <= SYNTHESIZED_WIRE_19;
Q6 <= SYNTHESIZED_WIRE_21;
Q7 <= SYNTHESIZED_WIRE_22;
SYNTHESIZED_WIRE_5 <= '0';
SYNTHESIZED_WIRE_24 <= '0';




b2v_inst1 : 74157_0
PORT MAP(A1 => P0,
		 B1 => SYNTHESIZED_WIRE_0,
		 SEL => SYNTHESIZED_WIRE_25,
		 B2 => SYNTHESIZED_WIRE_2,
		 A3 => P2,
		 B3 => SYNTHESIZED_WIRE_26,
		 A2 => P1,
		 B4 => SYNTHESIZED_WIRE_4,
		 GN => SYNTHESIZED_WIRE_5,
		 A4 => P3,
		 Y2 => SYNTHESIZED_WIRE_9,
		 Y1 => SYNTHESIZED_WIRE_10,
		 Y4 => SYNTHESIZED_WIRE_11,
		 Y3 => SYNTHESIZED_WIRE_8);


SYNTHESIZED_WIRE_27 <= NOT(SYNTHESIZED_WIRE_6);



b2v_inst2 : 74195_1
PORT MAP(ST/LDN => SYNTHESIZED_WIRE_27,
		 KN => SERIAL,
		 CLRN => MR,
		 D2 => SYNTHESIZED_WIRE_8,
		 D1 => SYNTHESIZED_WIRE_9,
		 D0 => SYNTHESIZED_WIRE_10,
		 J => SERIAL,
		 CLK => clock,
		 D3 => SYNTHESIZED_WIRE_11,
		 Q3 => SYNTHESIZED_WIRE_26,
		 Q0 => SYNTHESIZED_WIRE_23,
		 Q1 => SYNTHESIZED_WIRE_0,
		 Q2 => SYNTHESIZED_WIRE_2);



SYNTHESIZED_WIRE_25 <= NOT(PSN);



b2v_inst4 : 74195_2
PORT MAP(ST/LDN => SYNTHESIZED_WIRE_27,
		 KN => SYNTHESIZED_WIRE_26,
		 CLRN => MR,
		 D2 => SYNTHESIZED_WIRE_14,
		 D1 => SYNTHESIZED_WIRE_15,
		 D0 => SYNTHESIZED_WIRE_16,
		 J => SYNTHESIZED_WIRE_26,
		 CLK => clock,
		 D3 => SYNTHESIZED_WIRE_18,
		 Q3 => SYNTHESIZED_WIRE_22,
		 Q0 => SYNTHESIZED_WIRE_4,
		 Q1 => SYNTHESIZED_WIRE_19,
		 Q2 => SYNTHESIZED_WIRE_21);


b2v_inst8 : 74157_3
PORT MAP(A1 => P4,
		 B1 => SYNTHESIZED_WIRE_19,
		 SEL => SYNTHESIZED_WIRE_25,
		 B2 => SYNTHESIZED_WIRE_21,
		 A3 => P6,
		 B3 => SYNTHESIZED_WIRE_22,
		 A2 => P5,
		 B4 => SYNTHESIZED_WIRE_23,
		 GN => SYNTHESIZED_WIRE_24,
		 A4 => P7,
		 Y2 => SYNTHESIZED_WIRE_15,
		 Y1 => SYNTHESIZED_WIRE_16,
		 Y4 => SYNTHESIZED_WIRE_18,
		 Y3 => SYNTHESIZED_WIRE_14);


SYNTHESIZED_WIRE_6 <= LRN OR PSN;


END bdf_type;